FirstChapter
0
easy
