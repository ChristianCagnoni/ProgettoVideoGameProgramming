FirstChapter
0
easy
lt
