FirstChapter
1
easy
